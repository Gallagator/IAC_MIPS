`include "package.v"

module mips_cpu_bus(
    /* Standard signals */
    input logic clk,
    input logic reset,
    output logic active,
    output logic[31:0] register_v0,

    /* Avalon memory mapped bus controller (master) */
    output logic[31:0] address,
    output logic write,
    output logic read,
    input logic waitrequest,
    output logic[31:0] writedata,
    output logic[3:0] byteenable,
    input logic[31:0] readdata
);
    /* readdata/writedata big endian */
    logic[31:0] readdata_eb;
    logic[31:0] writedata_eb;

    /* Program Counter, instruction register, state */
    logic[31: 0] pc, pc_branch;
    branch_delay_state_t branch_delayed;

    logic[31: 0] ir, effective_ir;
    state_t state;

    /* Register file outputs */  
    logic[31:0] rs_val, rt_val;

    /* Reg file inputs */
    logic reg_file_write;
    logic[31:0] reg_file_data_in;
    logic[4:0] reg_file_rs;
    logic[4:0] reg_file_rt;
    logic[4:0] reg_file_rd;

    /* ALU */
    logic[31:0] alu_out;
    logic[5:0] alu_fncode;
    logic[31:0] alu_a;
    logic[31:0] alu_b;

    /* Instruction decode */
    logic[2:0] instr_type;
    logic[5:0] opcode;

    /* rtype instructions */
    logic[4:0] rtype_rs;
    logic[4:0] rtype_rt;
    logic[4:0] rtype_rd;
    logic[4:0] rtype_shamnt;
    logic[31:0] extended_shamnt;
    logic immediate_shift;
    logic[5:0] rtype_fncode;
    

    /* itype instructions */
    logic[4:0] itype_rs;
    logic[4:0] itype_rt;
    logic[31:0] itype_immediate;
    logic[31:0] loadstore_word; // bytes_control output.
    logic[3:0] bytes_byteenable;    // bytes_control output.

    /* jtype_instructions */
    logic[25:0] jtype_address;

    logic waitrequest_prev;

    assign opcode = effective_ir[31:26];

    /* rtype */
    assign rtype_rs     = effective_ir[25:21];
    assign rtype_rt     = effective_ir[20:16];
    assign rtype_rd     = effective_ir[15:11];
    assign rtype_shamnt = effective_ir[10:6];
    assign extended_shamnt = {27'b0, rtype_shamnt};
    assign rtype_fncode = effective_ir[5:0];

    /* itype */
    assign itype_rs     = effective_ir[25:21];
    assign itype_rt     = effective_ir[20:16];

    /* jtype */
    assign jtype_address = effective_ir[25:0];

    /* Bit addressing does not work in  always comb blocks. */
    always_comb begin
        
        /* Set active signal. pc must not be 0 and instruction must not 
         * have finished. */
        active = pc != 0 || state != STATE_FETCH;
        /* Decoding */
        /* Grabs the instruction that has just been fetched. */
        effective_ir = (state == STATE_EXECUTE && !waitrequest_prev) 
                       ? readdata_eb : ir;

        if(opcode == OPCODE_RTYPE) begin 
            immediate_shift = rtype_fncode == FUNCT_SLL || 
                              rtype_fncode == FUNCT_SRL || 
                              rtype_fncode == FUNCT_SRA;

            instr_type = RTYPE;
            reg_file_rs = rtype_rs;
            reg_file_rt = rtype_rt;
            reg_file_rd = rtype_rd;
            reg_file_write = state == STATE_EXECUTE;
            reg_file_data_in = alu_out;
            alu_a = immediate_shift ? extended_shamnt : rs_val;
            alu_b = rt_val;
        end
        else if(opcode == OPCODE_J || opcode == OPCODE_JAL) begin
            instr_type = JTYPE;
        end
        else begin
            instr_type = ITYPE;
            reg_file_rs = itype_rs;
            reg_file_rt = itype_rt;  // Mysteriously needed.
            reg_file_rd = itype_rt;

            if(reg_file_rt == 5'b10001) begin
                reg_file_rd = 31;
            end

            alu_a = rs_val;
            alu_b = itype_immediate;
        end

        case(state) 
            STATE_FETCH: begin
                reg_file_write = 0;
                read = 1;
                write = 0;
                address = pc;
                byteenable = 4'b1111;
            end
            STATE_EXECUTE : begin

                if(opcode == OPCODE_BEQ || opcode == OPCODE_BGTZ || opcode == OPCODE_BLEZ) begin
                    alu_a = itype_immediate;
                    alu_b = pc;
                    $display("CPU   alu_a: %x, alu_b: %x", alu_a, alu_b);
                end

                else if(opcode == OPCODE_REGIMM) begin
                    alu_a = itype_immediate;
                    alu_b = pc;
                    //$display("CPU   reg_file_rt: %b", reg_file_rt);
                    if(reg_file_rt == 5'b10001 || reg_file_rt == 5'b10000) begin   // BGEZAL and BLTZAL
                        reg_file_write = 1;
                        reg_file_data_in = pc+4;
                        $display("CPU   reg_file_data_in: %x", reg_file_data_in);
                    end

                end


                else if(opcode == OPCODE_LW) begin
                    write = 0;
                    read = 1;
                    byteenable = 4'b1111;
                    address = alu_out;
                    reg_file_write = 0;
                end
                
                else if(opcode == OPCODE_SW) begin
                    write = 0; 
                    read = 0;
                    byteenable = 4'b1111;
                    address = alu_out;
                    writedata_eb = rt_val;
                    reg_file_write = 0;
                end
                else if(opcode == OPCODE_LBU || opcode == OPCODE_LB || 
                        opcode == OPCODE_LHU || opcode == OPCODE_LH || 
                        opcode == OPCODE_LWL || opcode == OPCODE_LWR) begin     // Don't know if I can shorten this by putting it as default.
                    write = 0;
                    read = 1;
                    address = alu_out;
                    reg_file_write = 0;
                    byteenable = bytes_byteenable;
                end
                else if(opcode == OPCODE_LUI) begin
                    write = 0;
                    read = 0;
                    reg_file_data_in = itype_immediate;
                    reg_file_write = 1;
                end
                else begin
                    write = 0;  
                    read = 0;
                    reg_file_write = 1;
                    reg_file_data_in = alu_out;
                end

            end
            STATE_MEMORY : begin
                reg_file_write = 1;
                case(opcode)
                    OPCODE_LW : begin
                        reg_file_data_in = readdata_eb;
                    end
                    OPCODE_SW : begin
                        write = 1;
                    end
                    default : begin     // LBU, LB, LHU, LH, LWL, LWR
                        reg_file_data_in = loadstore_word;
                    end
                endcase
            end
        endcase

    end

    always @(state) begin
        case(state)
            STATE_FETCH : $display("-----------------------------------------\nSTATE FETCH");
            STATE_EXECUTE : $display("STATE EXECUTE");
            STATE_MEMORY : $display("STATE MEMORY");
        endcase
    end

    always @(pc) begin
        $display("CPU   pc: %x", pc);
    end

    always @(posedge clk) begin
        waitrequest_prev <= waitrequest;
       
        if(reset) begin
            pc <= 32'hBFC0_0000;
            state <= STATE_FETCH;
            pc_branch <= 0;
            branch_delayed <= BRANCH_NONE;
        end
        else if(active) begin
            case(state)  
                STATE_FETCH : begin
                    //reg_file_write <= 0;
                    /* Won't exit the fetch state if bus isn't ready to be
                     * read from yet. Further, it won't do anything if 
                     * it's still waiting */ 
                    if(!waitrequest) begin
                        pc <= pc + 4;
                        state <= STATE_EXECUTE;
                    end

                end
                STATE_EXECUTE : begin
                    ir <= waitrequest_prev ? ir : readdata_eb;

                    case(instr_type) 
                        RTYPE : begin
                            if(rtype_fncode == FUNCT_JR && branch_delayed == BRANCH_NONE) begin
                                pc_branch <= rs_val;
                                $display("JR");
                                $display("CPU   pc_branch: %x", pc_branch);
                                branch_delayed <= BRANCH_DELAYED;
                            end
                            state <= STATE_FETCH;
                        end 
                        ITYPE : begin

                            if(opcode == OPCODE_BEQ && rs_val == rt_val && branch_delayed == BRANCH_NONE) begin  // Else we go to Fetch state only.
                                pc_branch <= alu_out;
                                branch_delayed <= BRANCH_DELAYED;
                                state <= STATE_FETCH;
                                $display("BEQ");
                            end

                            else if(opcode == OPCODE_REGIMM) begin
                                 && $signed(rs_val) >= 0 && branch_delayed == BRANCH_NONE
                                if(reg_file_rt == 5'b00001 || reg_file_rt == 5'b10001 && $signed(rs_val) >= 0 && branch_delayed == BRANCH_NONE) begin   // BGEZ and BGEZAL
                                    pc_branch <= alu_out;
                                    branch_delayed <= BRANCH_DELAYED;
                                    
                                end
                    
                                else if(reg_file_rt == 5'b0 || reg_file_rt == 5'b10000 && $signed(rs_val) < 0 && branch_delayed == BRANCH_NONE) begin  // BLTZ
                                    pc_branch <= alu_out;
                                    branch_delayed <= BRANCH_DELAYED;
                                    
                                end 
                                
                                state <= STATE_FETCH;
                                $display("BGEZAL");
                                $display("CPU   alu_out: %x", alu_out);
                                $display("CPU   rs: %x", rs_val);
                            end
                            else if(opcode == OPCODE_BGTZ && $signed(rs_val) > 0 && branch_delayed == BRANCH_NONE) begin
                                pc_branch <= alu_out;
                                branch_delayed <= BRANCH_DELAYED;
                                $display("BGTZ");
                                $display("CPU   alu_out: %x", alu_out);
                                $display("CPU   rs: %x", rs_val);
                                state <= STATE_FETCH;

                            end

                            else if(opcode == OPCODE_BLEZ && $signed(rs_val) <= 0 && branch_delayed == BRANCH_NONE) begin
                                pc_branch <= alu_out;
                                branch_delayed <= BRANCH_DELAYED;
                                $display("BLEZ");
                                $display("CPU   alu_out: %x", alu_out);
                                $display("CPU   rs: %x", rs_val);
                                state <= STATE_FETCH;

                            end

                            /* Will also have to include other load instrs */
                            else if( opcode == OPCODE_LW || opcode == OPCODE_LBU || 
                                opcode == OPCODE_LB || opcode == OPCODE_LH || 
                                opcode == OPCODE_LHU || opcode == OPCODE_LWL || 
                                opcode == OPCODE_LWR ) begin    // Don't know I could make this shorter by putting it into the else statement.
                                
                                if(!waitrequest) begin
                                    state <= STATE_MEMORY;
                                end 
                            end
                            else if(opcode == OPCODE_SW) begin
                                if(!waitrequest) begin 
                                    state <= STATE_MEMORY;
                                end
                            end 
                            else begin
                                $display("ADDIU");
                                state <= STATE_FETCH;
                            end

                        end 
                        JTYPE : begin

                        end 
                        default : ;
                    endcase

                    if(branch_delayed == BRANCH_DELAYED) begin
                        pc <= pc_branch;
                        $display("BRANCH   pc: %x", pc);
                        branch_delayed <= BRANCH_NONE;
                    end
                    
                end
                STATE_MEMORY : begin
                    state <= STATE_FETCH;
                end

                default : ;
            endcase
        end
    end

    alu_ctrl alu_ctrl(.opcode(opcode),
                      .rtype_fncode(rtype_fncode),
                      .fncode(alu_fncode)
    );

    reg_file reg_file(.clk(clk), 
                      .reset(reset), 
                      .addr_a(reg_file_rs),
                      .addr_b(reg_file_rt),
                      .write_addr(reg_file_rd),
                      .write(reg_file_write),
                      .data_in(reg_file_data_in),
                      .a(rs_val),
                      .b(rt_val),
                      .register_v0(register_v0)
    );

    alu alu(.a(alu_a), .b(alu_b), .fncode(alu_fncode), .r(alu_out));

    toggle_endianness to_big(.a(readdata), .r(readdata_eb));
    toggle_endianness to_little(.a(writedata_eb), .r(writedata));

    sign_extension sign_extension(
        .itype_immediate(effective_ir[15:0]),
        .opcode(opcode),
        .signed_itype_immediate(itype_immediate)
    );

    bytes_control bytes_control(
        .readdata_eb(readdata_eb),
        .opcode(opcode),
        .lsb_bits(address[1:0]),
        .bytes_out(loadstore_word),
        .rt_val_itype(rt_val),
        .byteenable(bytes_byteenable)
    );

endmodule

module toggle_endianness(
    input logic[31:0] a,
    output logic[31:0] r
);
    assign r = {a[7:0], a[15:8], a[23:16], a[31:24]};
 
endmodule
