module alu_control(
    input logic[1:0] aluop,
    input logic[4:0] funct,
    output logic[3:0] op
);


    
endmodule